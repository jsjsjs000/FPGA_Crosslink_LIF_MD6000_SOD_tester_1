/*
This demo is for the CrossLink LIF-MD6000 on Lattice Semiconductor Master Link Board.
*/
module gpio_test(pin,reset);

output reg [3:0] pin;	//LEDs
input reset;			// Reset switch
//reg reset = 1; 

wire clk_osc;		// Signal from internal oscillator i.e 6 MHz
reg [25:0] clk_f = 0;	//count Register to achieve  i.e 2.86 Hz which is visible to human eyes

//------------------------- Internal Oscillator----------------------------------
/*	OSCI runs at 10 KHz in low frequency mode and at maximum 48 MHz in high frequency mode with output divider by 1, 2, 4 or 8.
	The HFCLKOUT will be 48/8 = 6 MHz (166.66 ns).
*/
defparam I1.HFCLKDIV = 1; // 1,2,4,8 - Divider value for HFCLKOUT signal. Output is divided by 8 here.
OSCI I1 (
.HFOUTEN(1'b1),			// Enable signal for HFCLKOUT. 
.HFCLKOUT(clk_osc),		// High frequency output. Used as the base clock for this demo
.LFCLKOUT(LFCLKOUT));	// Low frequency output. Not used in this demo
//--------------------------------------------------------------------------------


//------------------------- Counter----------------------------------
/* 	A counter is used to slow down the clock for LED shifting logic.
	This actually works as a clock divider with a larger value.
	This is needed because the toggling of an LED at 6 MHz (166.66 ns) cannot be seen by human eyes.
*/
always @ (posedge clk_osc)
	begin
		clk_f<=clk_f+1'b1;	// Counter
	end
//-------------------------------------------------------------------



//------------------------- Shift register ---------------------------
/*
	A walking 1s pattern is generated by shifting "1101" left in each clock cycle.
	A synchronous reset is used to bring back the LEDs to initial state.
	The clock to this logic is the 20th bit of the counter register.
	The clock to this logic is a slower clock made using a counter.
*/
	always @ (posedge clk_f[20])
		begin
			if (reset==0)
				pin<=4'b1110; //"1001"; 		// Initial value of LEDs.
			else 
				pin<={pin[0],pin[3:1]}; // Shifting the LED values to make a walking 1s pattern
		end	
//-------------------------------------------------------------------
endmodule